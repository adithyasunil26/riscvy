module execute(
  input [63:0] a,
  input [63:0] readdata1,
  input [63:0] readdata2,
);

endmodule